library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library work;
use work.riscv_pkg.all;

entity execute is
    Port (
        -- Inputs
	i_clk 	      : in std_logic;
i_alu_op      : in  std_logic_vector(2 downto 0);
        i_rs1_data    : in  STD_LOGIC_VECTOR(31 downto 0);
        i_rs2_data    : in  STD_LOGIC_VECTOR(31 downto 0);
        i_imm         : in  STD_LOGIC_VECTOR(31 downto 0);
        i_pc          : in  STD_LOGIC_VECTOR(31 downto 0);
        i_src_imm     : in  STD_LOGIC;
        i_branch      : in  STD_LOGIC;
        i_jump        : in  STD_LOGIC;
	




        -- Outputs
        o_pc_transfer : out STD_LOGIC_VECTOR(31 downto 0);
        o_alu_result  : out STD_LOGIC_VECTOR(31 downto 0);
        o_store_data  : out STD_LOGIC_VECTOR(31 downto 0);
        o_pc_target   : out STD_LOGIC_VECTOR(31 downto 0)
    );
end execute;

architecture Behavioral of execute is


component riscv_adder is
  generic (
    N : positive := 32
  );
  port (
    i_a    : in  std_logic_vector(N-1 downto 0);
    i_b    : in  std_logic_vector(N-1 downto 0);
    i_sign : in  std_logic;
    i_sub  : in  std_logic;
    o_sum  : out std_logic_vector(N downto 0)
 
  );
end component riscv_adder;

component riscv_alu is
  port (
    i_arith  : in  std_logic;                                -- Arith/Logic
    i_sign   : in  std_logic;                                -- Signed/Unsigned
    i_opcode : in  std_logic_vector(2 downto 0); -- ALU opcodes
    i_shamt  : in  std_logic_vector(SHAMT_WIDTH-1 downto 0); -- Shift Amount
    i_src1   : in  std_logic_vector(XLEN-1 downto 0);        -- Operand A
    i_src2   : in  std_logic_vector(XLEN-1 downto 0);        -- Operand B
    o_res    : out std_logic_vector(XLEN-1 downto 0));       -- Result
end component riscv_alu;


    -- Intermediate signals
    signal alu_in2      : STD_LOGIC_VECTOR(31 downto 0);
    signal alu_out      : STD_LOGIC_VECTOR(31 downto 0);
    signal adder_out    : STD_LOGIC_VECTOR(32 downto 0);  -- Result of the adder
    signal pc_target    : STD_LOGIC_VECTOR(31 downto 0);
    
begin
    -- **S�lection entre rs2_data et imm pour l'ALU (src_imm)**
    alu_in2 <= i_imm when i_src_imm = '1' else i_rs2_data;

    -- ALU instance
    ALU_INST : riscv_alu
        port map (
            i_arith  => '1', -- Assuming arithmetic operation
            i_sign   => '1', -- Assuming signed operation
            i_opcode => i_alu_op,
            i_shamt  => i_imm(4 downto 0), -- Extract shift amount
            i_src1   => i_rs1_data,
            i_src2   => alu_in2,
            o_res    => alu_out
        );

    -- **Adder instance for PC target calculation**
    ADDER_INST : riscv_adder
        generic map (
            N => 32
        )
        port map (
            i_a    => i_pc,
            i_b    => i_imm,
            i_sign => '1',     -- Assuming signed addition
            i_sub  => '0',     -- No subtraction
            o_sum  => adder_out
        );

process(i_clk)
begin
if rising_edge(i_clk) then
    o_alu_result <= alu_out;
    o_store_data <= i_rs2_data;
end if;
end process;
    o_pc_target  <= adder_out(31 downto 0); -- Discard the carry bit
    o_pc_transfer <= adder_out(31 downto 0) when (i_jump = '1' or i_branch = '1') else alu_out;
o_pc_transfer <= alu_out when (i_jump = '1' or i_branch = '1')else (i_pc + 4);

end Behavioral;
